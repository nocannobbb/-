`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2018/12/06 17:05:04
// Design Name: 
// Module Name: floprc
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


//floprc #(5) r4E(clk,rst,flushE,rsD,rsE);

module floprc #(parameter WIDTH = 8)(
	input wire clk,rst,flush,
	input wire [WIDTH-1:0] d,
	output reg [WIDTH-1:0] q
    );

	always @(posedge clk or posedge rst) begin
		if(rst) begin
			q <= 0;
		end

		else if(flush) begin
			q <= 0;
		end

		else begin
			q <= d;
		end
	end
endmodule
